�� 
 m o d u l e   m e m   # (                                       / /    
         p a r a m e t e r     A D D R _ L E N     =   1 1       / /    
 )   (  
         i n p u t     c l k ,   r s t ,  
         i n p u t     [ A D D R _ L E N - 1 : 0 ]   a d d r ,   / /   m e m o r y   a d d r e s s  
         o u t p u t   r e g   [ 3 1 : 0 ]   r d _ d a t a ,     / /   d a t a   r e a d   o u t  
         i n p u t     w r _ r e q ,  
         i n p u t     [ 3 1 : 0 ]   w r _ d a t a               / /   d a t a   w r i t e   i n  
 ) ;  
 l o c a l p a r a m   M E M _ S I Z E   =   1 < < A D D R _ L E N ;  
 r e g   [ 3 1 : 0 ]   r a m _ c e l l   [ M E M _ S I Z E ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k   o r   p o s e d g e   r s t )  
         i f ( r s t )  
                 r d _ d a t a   < =   0 ;  
         e l s e  
                 r d _ d a t a   < =   r a m _ c e l l [ a d d r ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k )  
         i f ( w r _ r e q )    
                 r a m _ c e l l [ a d d r ]   < =   w r _ d a t a ;  
  
 i n i t i a l   b e g i n  
         / /   d s t   m a t r i x   C  
         r a m _ c e l l [               0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 9 2 1 b 2 3 6 ;  
         r a m _ c e l l [               1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 6 f 9 2 d f 6 ;  
         r a m _ c e l l [               2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 3 9 a 3 9 6 8 ;  
         r a m _ c e l l [               3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 3 5 c 7 4 b b ;  
         r a m _ c e l l [               4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 3 7 a 6 d d 8 ;  
         r a m _ c e l l [               5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 3 8 a c 5 c 6 ;  
         r a m _ c e l l [               6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 2 f d 5 8 8 9 ;  
         r a m _ c e l l [               7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f f 9 e 5 6 d 7 ;  
         r a m _ c e l l [               8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 d 0 f 9 6 5 a ;  
         r a m _ c e l l [               9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 5 3 7 1 9 0 a ;  
         r a m _ c e l l [             1 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b c 6 a 0 4 c 6 ;  
         r a m _ c e l l [             1 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 2 c 8 3 e 4 4 ;  
         r a m _ c e l l [             1 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 3 8 a a e 5 1 ;  
         r a m _ c e l l [             1 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 5 9 1 9 c 6 e ;  
         r a m _ c e l l [             1 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 7 7 c 7 5 5 f ;  
         r a m _ c e l l [             1 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 f 6 b 6 c b e ;  
         r a m _ c e l l [             1 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 6 3 6 7 9 e 5 ;  
         r a m _ c e l l [             1 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 4 b b 6 b 7 e ;  
         r a m _ c e l l [             1 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 2 7 d 9 a 9 3 ;  
         r a m _ c e l l [             1 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 2 1 1 7 d 2 7 ;  
         r a m _ c e l l [             2 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 b 6 a 7 b e 2 ;  
         r a m _ c e l l [             2 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 2 c e b c 8 5 ;  
         r a m _ c e l l [             2 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f c a 8 f f 8 a ;  
         r a m _ c e l l [             2 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 3 d 3 b 2 5 c ;  
         r a m _ c e l l [             2 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 f 1 2 1 c 4 a ;  
         r a m _ c e l l [             2 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 4 6 d 8 4 3 b ;  
         r a m _ c e l l [             2 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 3 2 c d a 3 7 ;  
         r a m _ c e l l [             2 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 a 8 8 1 c 2 d ;  
         r a m _ c e l l [             2 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 5 6 b c 2 d a ;  
         r a m _ c e l l [             2 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 a 4 f a b b b ;  
         r a m _ c e l l [             3 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 4 8 2 8 3 9 9 ;  
         r a m _ c e l l [             3 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 1 9 6 9 b 2 1 ;  
         r a m _ c e l l [             3 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 c 2 1 5 d 9 3 ;  
         r a m _ c e l l [             3 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 5 0 b c 6 5 d ;  
         r a m _ c e l l [             3 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 4 d f 6 c 7 4 ;  
         r a m _ c e l l [             3 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 5 1 9 a 6 1 8 ;  
         r a m _ c e l l [             3 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 1 9 5 8 0 9 b ;  
         r a m _ c e l l [             3 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 7 d 6 5 4 b d ;  
         r a m _ c e l l [             3 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 6 d b f a 7 7 ;  
         r a m _ c e l l [             3 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e a 6 5 5 8 f 7 ;  
         r a m _ c e l l [             4 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 1 d b 0 0 8 2 ;  
         r a m _ c e l l [             4 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 c 4 5 8 7 5 5 ;  
         r a m _ c e l l [             4 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 0 5 6 0 d 3 8 ;  
         r a m _ c e l l [             4 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 8 0 1 6 7 f b ;  
         r a m _ c e l l [             4 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 7 c 4 4 3 5 5 ;  
         r a m _ c e l l [             4 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 a d 6 1 6 6 4 ;  
         r a m _ c e l l [             4 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 c 0 3 e 5 a a ;  
         r a m _ c e l l [             4 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c c 9 1 3 3 1 f ;  
         r a m _ c e l l [             4 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 c 4 6 3 3 2 f ;  
         r a m _ c e l l [             4 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 4 4 c 1 0 1 4 ;  
         r a m _ c e l l [             5 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 7 5 4 a c f 8 ;  
         r a m _ c e l l [             5 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 b 5 0 d e 2 6 ;  
         r a m _ c e l l [             5 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 7 4 d c 1 0 3 ;  
         r a m _ c e l l [             5 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 0 c 3 e 7 c 8 ;  
         r a m _ c e l l [             5 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a e 3 e 7 c c 3 ;  
         r a m _ c e l l [             5 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 2 7 0 5 7 c 3 ;  
         r a m _ c e l l [             5 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 0 2 0 0 2 4 7 ;  
         r a m _ c e l l [             5 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 9 e b 0 9 3 8 ;  
         r a m _ c e l l [             5 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 7 4 1 2 d 8 b ;  
         r a m _ c e l l [             5 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 f c 1 1 5 7 1 ;  
         r a m _ c e l l [             6 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 0 2 8 9 2 a e ;  
         r a m _ c e l l [             6 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d e f 7 8 a 3 f ;  
         r a m _ c e l l [             6 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 0 b a 6 2 5 a ;  
         r a m _ c e l l [             6 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 4 4 b a 7 0 c ;  
         / /   s r c   m a t r i x   A  
         r a m _ c e l l [             6 4 ]   =   3 2 ' h 4 1 7 c 8 b 8 9 ;  
         r a m _ c e l l [             6 5 ]   =   3 2 ' h 8 8 d a a c 7 8 ;  
         r a m _ c e l l [             6 6 ]   =   3 2 ' h 9 a 2 4 b f 4 9 ;  
         r a m _ c e l l [             6 7 ]   =   3 2 ' h d 4 2 3 6 f 6 4 ;  
         r a m _ c e l l [             6 8 ]   =   3 2 ' h 0 d 9 3 9 6 b e ;  
         r a m _ c e l l [             6 9 ]   =   3 2 ' h 8 4 7 d 3 3 d f ;  
         r a m _ c e l l [             7 0 ]   =   3 2 ' h c a b 4 a f 0 0 ;  
         r a m _ c e l l [             7 1 ]   =   3 2 ' h b 4 1 c b 7 f 9 ;  
         r a m _ c e l l [             7 2 ]   =   3 2 ' h 9 1 1 d f b c 2 ;  
         r a m _ c e l l [             7 3 ]   =   3 2 ' h 1 9 d 5 a 0 e a ;  
         r a m _ c e l l [             7 4 ]   =   3 2 ' h 6 d 5 b 4 7 e 6 ;  
         r a m _ c e l l [             7 5 ]   =   3 2 ' h d 2 a 5 b f 6 d ;  
         r a m _ c e l l [             7 6 ]   =   3 2 ' h f f 2 f e 5 c c ;  
         r a m _ c e l l [             7 7 ]   =   3 2 ' h 6 4 5 b 9 b 6 c ;  
         r a m _ c e l l [             7 8 ]   =   3 2 ' h b a 7 e 5 7 3 9 ;  
         r a m _ c e l l [             7 9 ]   =   3 2 ' h c 3 5 9 9 5 6 b ;  
         r a m _ c e l l [             8 0 ]   =   3 2 ' h d 3 d 3 0 d 3 c ;  
         r a m _ c e l l [             8 1 ]   =   3 2 ' h 0 1 4 d 6 4 c e ;  
         r a m _ c e l l [             8 2 ]   =   3 2 ' h 1 6 4 5 e b 3 6 ;  
         r a m _ c e l l [             8 3 ]   =   3 2 ' h d 0 c 6 6 4 7 7 ;  
         r a m _ c e l l [             8 4 ]   =   3 2 ' h 6 d e 9 a 9 3 d ;  
         r a m _ c e l l [             8 5 ]   =   3 2 ' h f 6 3 9 3 9 0 a ;  
         r a m _ c e l l [             8 6 ]   =   3 2 ' h d 1 b 2 2 c 4 0 ;  
         r a m _ c e l l [             8 7 ]   =   3 2 ' h 1 4 d 1 b d 4 6 ;  
         r a m _ c e l l [             8 8 ]   =   3 2 ' h d 7 1 9 0 9 8 1 ;  
         r a m _ c e l l [             8 9 ]   =   3 2 ' h 0 e 6 4 b 2 e 6 ;  
         r a m _ c e l l [             9 0 ]   =   3 2 ' h 8 7 8 c e 5 8 4 ;  
         r a m _ c e l l [             9 1 ]   =   3 2 ' h 8 2 7 6 7 a e 8 ;  
         r a m _ c e l l [             9 2 ]   =   3 2 ' h 9 0 b 5 b d e 6 ;  
         r a m _ c e l l [             9 3 ]   =   3 2 ' h c 9 c 9 d 8 5 e ;  
         r a m _ c e l l [             9 4 ]   =   3 2 ' h c 6 7 a b c 5 2 ;  
         r a m _ c e l l [             9 5 ]   =   3 2 ' h b 0 1 e 8 9 0 3 ;  
         r a m _ c e l l [             9 6 ]   =   3 2 ' h f a 4 e 7 4 d 5 ;  
         r a m _ c e l l [             9 7 ]   =   3 2 ' h 3 3 e 0 9 f b f ;  
         r a m _ c e l l [             9 8 ]   =   3 2 ' h 5 f 1 c 3 c 6 4 ;  
         r a m _ c e l l [             9 9 ]   =   3 2 ' h c 1 a e 3 5 e b ;  
         r a m _ c e l l [           1 0 0 ]   =   3 2 ' h 2 2 c 5 d 5 1 9 ;  
         r a m _ c e l l [           1 0 1 ]   =   3 2 ' h c f 4 6 4 6 4 f ;  
         r a m _ c e l l [           1 0 2 ]   =   3 2 ' h 5 b c 4 1 6 a e ;  
         r a m _ c e l l [           1 0 3 ]   =   3 2 ' h 0 7 e 7 d b 3 1 ;  
         r a m _ c e l l [           1 0 4 ]   =   3 2 ' h a 7 8 6 8 6 a 0 ;  
         r a m _ c e l l [           1 0 5 ]   =   3 2 ' h e f d e 0 1 0 b ;  
         r a m _ c e l l [           1 0 6 ]   =   3 2 ' h a 6 2 9 e a 6 8 ;  
         r a m _ c e l l [           1 0 7 ]   =   3 2 ' h 3 7 1 3 0 d 1 c ;  
         r a m _ c e l l [           1 0 8 ]   =   3 2 ' h e b 5 9 f c 2 9 ;  
         r a m _ c e l l [           1 0 9 ]   =   3 2 ' h b a 3 9 2 6 c 2 ;  
         r a m _ c e l l [           1 1 0 ]   =   3 2 ' h 6 a 2 0 f 3 4 0 ;  
         r a m _ c e l l [           1 1 1 ]   =   3 2 ' h 3 f 5 a b f 0 a ;  
         r a m _ c e l l [           1 1 2 ]   =   3 2 ' h e b 6 b 1 e a 4 ;  
         r a m _ c e l l [           1 1 3 ]   =   3 2 ' h 1 a 3 2 7 0 c 9 ;  
         r a m _ c e l l [           1 1 4 ]   =   3 2 ' h 9 b c d 4 b 8 2 ;  
         r a m _ c e l l [           1 1 5 ]   =   3 2 ' h c 1 5 f 2 a c 1 ;  
         r a m _ c e l l [           1 1 6 ]   =   3 2 ' h 8 b a 3 2 7 4 7 ;  
         r a m _ c e l l [           1 1 7 ]   =   3 2 ' h 8 e 0 d 8 7 0 6 ;  
         r a m _ c e l l [           1 1 8 ]   =   3 2 ' h d 3 2 2 1 d 7 1 ;  
         r a m _ c e l l [           1 1 9 ]   =   3 2 ' h 5 9 8 7 8 1 5 c ;  
         r a m _ c e l l [           1 2 0 ]   =   3 2 ' h f b 3 0 0 e 4 5 ;  
         r a m _ c e l l [           1 2 1 ]   =   3 2 ' h 8 3 3 8 a a 4 a ;  
         r a m _ c e l l [           1 2 2 ]   =   3 2 ' h 9 7 f a f 7 b e ;  
         r a m _ c e l l [           1 2 3 ]   =   3 2 ' h 7 b 3 d 8 2 e c ;  
         r a m _ c e l l [           1 2 4 ]   =   3 2 ' h 3 d d 4 5 2 9 d ;  
         r a m _ c e l l [           1 2 5 ]   =   3 2 ' h 8 2 a 3 f 4 8 8 ;  
         r a m _ c e l l [           1 2 6 ]   =   3 2 ' h 2 4 1 f d 8 0 8 ;  
         r a m _ c e l l [           1 2 7 ]   =   3 2 ' h 6 0 f d 1 8 a a ;  
         / /   s r c   m a t r i x   B  
         r a m _ c e l l [           1 2 8 ]   =   3 2 ' h 3 1 0 3 1 f 0 f ;  
         r a m _ c e l l [           1 2 9 ]   =   3 2 ' h 8 0 2 0 9 5 3 0 ;  
         r a m _ c e l l [           1 3 0 ]   =   3 2 ' h 2 6 a 1 c 7 9 f ;  
         r a m _ c e l l [           1 3 1 ]   =   3 2 ' h 9 f 2 f 6 3 2 2 ;  
         r a m _ c e l l [           1 3 2 ]   =   3 2 ' h f 9 e b 4 1 3 f ;  
         r a m _ c e l l [           1 3 3 ]   =   3 2 ' h 8 1 d 6 f b e 7 ;  
         r a m _ c e l l [           1 3 4 ]   =   3 2 ' h 5 3 6 3 8 5 0 3 ;  
         r a m _ c e l l [           1 3 5 ]   =   3 2 ' h 4 b c 2 3 f d b ;  
         r a m _ c e l l [           1 3 6 ]   =   3 2 ' h 5 8 4 d c d 2 e ;  
         r a m _ c e l l [           1 3 7 ]   =   3 2 ' h f a 8 b 8 4 b 9 ;  
         r a m _ c e l l [           1 3 8 ]   =   3 2 ' h 2 f 3 0 d f d 4 ;  
         r a m _ c e l l [           1 3 9 ]   =   3 2 ' h 5 0 5 e c e 0 4 ;  
         r a m _ c e l l [           1 4 0 ]   =   3 2 ' h 7 2 6 8 c 4 4 e ;  
         r a m _ c e l l [           1 4 1 ]   =   3 2 ' h 0 e a a 9 a c a ;  
         r a m _ c e l l [           1 4 2 ]   =   3 2 ' h 1 4 9 6 3 c d b ;  
         r a m _ c e l l [           1 4 3 ]   =   3 2 ' h 1 6 6 b 1 4 8 6 ;  
         r a m _ c e l l [           1 4 4 ]   =   3 2 ' h d d f 0 b f 3 2 ;  
         r a m _ c e l l [           1 4 5 ]   =   3 2 ' h 1 3 d f 6 3 2 6 ;  
         r a m _ c e l l [           1 4 6 ]   =   3 2 ' h 7 d a 8 d e 7 d ;  
         r a m _ c e l l [           1 4 7 ]   =   3 2 ' h 0 9 c b c e 1 6 ;  
         r a m _ c e l l [           1 4 8 ]   =   3 2 ' h b 0 b 2 7 0 c 5 ;  
         r a m _ c e l l [           1 4 9 ]   =   3 2 ' h 8 a 4 2 0 2 d 2 ;  
         r a m _ c e l l [           1 5 0 ]   =   3 2 ' h c 1 e 2 2 0 d 7 ;  
         r a m _ c e l l [           1 5 1 ]   =   3 2 ' h 1 4 e b 5 a 4 2 ;  
         r a m _ c e l l [           1 5 2 ]   =   3 2 ' h f 9 f 5 3 4 c d ;  
         r a m _ c e l l [           1 5 3 ]   =   3 2 ' h 3 7 f 8 f 2 c 8 ;  
         r a m _ c e l l [           1 5 4 ]   =   3 2 ' h 5 3 e e 1 4 6 7 ;  
         r a m _ c e l l [           1 5 5 ]   =   3 2 ' h d d 9 c 2 d 5 2 ;  
         r a m _ c e l l [           1 5 6 ]   =   3 2 ' h e 4 3 c 5 7 2 1 ;  
         r a m _ c e l l [           1 5 7 ]   =   3 2 ' h 0 b 3 1 6 2 9 b ;  
         r a m _ c e l l [           1 5 8 ]   =   3 2 ' h 0 2 7 c 8 4 c f ;  
         r a m _ c e l l [           1 5 9 ]   =   3 2 ' h f f 3 a 6 b 2 b ;  
         r a m _ c e l l [           1 6 0 ]   =   3 2 ' h 1 a b e 2 4 1 2 ;  
         r a m _ c e l l [           1 6 1 ]   =   3 2 ' h 0 c 4 d 9 b 5 2 ;  
         r a m _ c e l l [           1 6 2 ]   =   3 2 ' h 9 4 7 9 0 3 5 4 ;  
         r a m _ c e l l [           1 6 3 ]   =   3 2 ' h 5 9 5 c e e 9 b ;  
         r a m _ c e l l [           1 6 4 ]   =   3 2 ' h 2 2 f d 3 b a 9 ;  
         r a m _ c e l l [           1 6 5 ]   =   3 2 ' h 4 b 5 5 0 8 2 4 ;  
         r a m _ c e l l [           1 6 6 ]   =   3 2 ' h d 8 b 9 e c 5 d ;  
         r a m _ c e l l [           1 6 7 ]   =   3 2 ' h 2 5 8 5 2 9 8 d ;  
         r a m _ c e l l [           1 6 8 ]   =   3 2 ' h f a e 9 b c 4 6 ;  
         r a m _ c e l l [           1 6 9 ]   =   3 2 ' h e 4 0 0 8 c e b ;  
         r a m _ c e l l [           1 7 0 ]   =   3 2 ' h e 4 f b 7 7 4 6 ;  
         r a m _ c e l l [           1 7 1 ]   =   3 2 ' h 1 5 0 6 8 3 9 0 ;  
         r a m _ c e l l [           1 7 2 ]   =   3 2 ' h 0 6 6 4 3 e e d ;  
         r a m _ c e l l [           1 7 3 ]   =   3 2 ' h 8 4 e 5 9 2 0 9 ;  
         r a m _ c e l l [           1 7 4 ]   =   3 2 ' h e 8 a 6 e 5 0 7 ;  
         r a m _ c e l l [           1 7 5 ]   =   3 2 ' h 5 0 a 2 3 e 1 a ;  
         r a m _ c e l l [           1 7 6 ]   =   3 2 ' h 1 e c 4 0 2 1 0 ;  
         r a m _ c e l l [           1 7 7 ]   =   3 2 ' h a d 5 2 0 f 6 d ;  
         r a m _ c e l l [           1 7 8 ]   =   3 2 ' h 3 f 9 f 6 1 2 f ;  
         r a m _ c e l l [           1 7 9 ]   =   3 2 ' h 7 8 f e 0 0 f 5 ;  
         r a m _ c e l l [           1 8 0 ]   =   3 2 ' h 4 9 c c 7 4 8 d ;  
         r a m _ c e l l [           1 8 1 ]   =   3 2 ' h f 7 1 2 5 5 c b ;  
         r a m _ c e l l [           1 8 2 ]   =   3 2 ' h a 8 5 3 7 d e c ;  
         r a m _ c e l l [           1 8 3 ]   =   3 2 ' h d 1 6 e 0 e 7 3 ;  
         r a m _ c e l l [           1 8 4 ]   =   3 2 ' h 9 5 b a 4 1 6 b ;  
         r a m _ c e l l [           1 8 5 ]   =   3 2 ' h 8 8 5 9 4 1 a 7 ;  
         r a m _ c e l l [           1 8 6 ]   =   3 2 ' h d 9 0 9 3 0 8 a ;  
         r a m _ c e l l [           1 8 7 ]   =   3 2 ' h 5 a 2 f e 0 5 3 ;  
         r a m _ c e l l [           1 8 8 ]   =   3 2 ' h d 3 f 1 4 f b 3 ;  
         r a m _ c e l l [           1 8 9 ]   =   3 2 ' h b 8 4 6 3 6 9 6 ;  
         r a m _ c e l l [           1 9 0 ]   =   3 2 ' h e a 2 5 b c 8 c ;  
         r a m _ c e l l [           1 9 1 ]   =   3 2 ' h 5 6 c d c 9 4 a ;  
 e n d  
  
 e n d m o d u l e  
  
 